module rca_pipe_2bit(a,b,cin,clk,sum,cout);
  input [7:0] a,b;
  input cin,clk;
  output [7:0] sum;
  output cout;


 endmodule
